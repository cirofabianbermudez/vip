`ifndef GPIO_UVC_SEQUENCER_SV
`define GPIO_UVC_SEQUENCER_SV

typedef uvm_sequencer #(gpio_uvc_sequence_item) gpio_uvc_sequencer;

`endif // GPIO_UVC_SEQUENCER_SV
