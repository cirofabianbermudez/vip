`ifndef I2C_UVC_SEQUENCER_SV
`define I2C_UVC_SEQUENCER_SV

typedef uvm_sequencer#(i2c_uvc_sequence_item) i2c_uvc_sequencer;

`endif  // I2C_UVC_SEQUENCER_SV
