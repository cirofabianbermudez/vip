`ifndef GPIO_UVC_CONFIG_SV
`define GPIO_UVC_CONFIG_SV

class gpio_uvc_config extends uvm_object;

  `uvm_object_utils(gpio_uvc_config)

  uvm_active_passive_enum  is_active = UVM_ACTIVE;
  bit                      coverage_enable;    

  extern function new(string name = "");

endclass : gpio_uvc_config

function gpio_uvc_config::new(string name = "");
  super.new(name);
endfunction : new

`endif // GPIO_UVC_CONFIG_SV
