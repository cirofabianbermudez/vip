`ifndef GPIO_UVC_MONITOR_SV
`define GPIO_UVC_MONITOR_SV

class gpio_uvc_monitor #(int WIDTH = 8) extends uvm_monitor;

  typedef gpio_uvc_monitor #(WIDTH) gpio_uvc_monitor_t;
  `uvm_component_param_utils(gpio_uvc_monitor_t)

  typedef virtual gpio_uvc_if #(WIDTH) gpio_uvc_if_t;
  gpio_uvc_if_t vif;

  uvm_analysis_port #(gpio_uvc_sequence_item) analysis_port;
  gpio_uvc_sequence_item trans;

  extern function new(string name, uvm_component parent);
  extern function void build_phase(uvm_phase phase);
  extern task run_phase(uvm_phase phase);
  extern task do_mon();

endclass : gpio_uvc_monitor


function gpio_uvc_monitor::new(string name, uvm_component parent);
  super.new(name, parent);
endfunction : new


function void gpio_uvc_monitor::build_phase(uvm_phase phase);
  if ( !uvm_config_db #(gpio_uvc_if_t)::get(get_parent(), "", "vif", vif) ) begin
		  `uvm_fatal(get_name(), "Could not retrieve gpio_uvc_if from config db")
	end

  analysis_port = new("analysis_port", this);

endfunction : build_phase


task gpio_uvc_monitor::run_phase(uvm_phase phase);
  trans = gpio_uvc_sequence_item::type_id::create("trans");
  do_mon();
endtask : run_phase


task gpio_uvc_monitor::do_mon();
  forever begin
    @(vif.gpio_pin)
    trans.gpio_pin = vif.gpio_pin;
    `uvm_info(get_type_name(), {"Got item ", trans.convert2string()}, UVM_MEDIUM)
    analysis_port.write(trans);
  end
endtask : do_mon

`endif // GPIO_UVC_MONITOR_SV
